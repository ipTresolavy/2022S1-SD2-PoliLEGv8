../Dataflow/shift_register.vhd