../ALU_4/ALU_4.vhd