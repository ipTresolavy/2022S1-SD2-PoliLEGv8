../Dataflow/data_memory_tb.vhd