../Dataflow/sign_extension_unit.vhd