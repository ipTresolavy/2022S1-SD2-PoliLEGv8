../Dataflow/ALU_pc.vhd