../Dataflow/sign_extension_unit_tb.vhd