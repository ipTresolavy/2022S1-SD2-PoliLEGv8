../ALU/ALU.vhd