../ALU/barrel_shifter_tb.vhd