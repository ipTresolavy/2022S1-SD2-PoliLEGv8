../ALU/PFA_tb.vhd