../Mul_Div_Unit/shift_register.vhd