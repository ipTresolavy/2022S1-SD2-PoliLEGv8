../ALU/ALU_tb.vhd