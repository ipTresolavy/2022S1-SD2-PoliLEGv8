../ALU/mul_div_unit.vhd