../ALU/mux4x1.vhd