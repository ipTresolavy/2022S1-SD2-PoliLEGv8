../ALU/alu.vhd