../Dataflow/instruction_memory_tb.vhd