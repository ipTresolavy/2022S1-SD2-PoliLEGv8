../Memory/instruction_memory_tb.vhd