../Dataflow/two_bit_left_shifter.vhd