../Control_Unit/control_unit.vhd