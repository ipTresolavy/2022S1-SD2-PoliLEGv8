../ALU/mux2x1_bin.vhd