../Dataflow/barrel_shifter.vhd