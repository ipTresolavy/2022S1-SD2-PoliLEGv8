../Dataflow/instruction_memory.vhd