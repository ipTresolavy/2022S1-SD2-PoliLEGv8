../Memory/data_memory.vhd