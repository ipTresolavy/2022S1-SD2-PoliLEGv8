../Two_Bit_Left_Shifter/two_bit_left_shifter.vhd