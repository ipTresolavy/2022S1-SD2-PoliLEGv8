../Dataflow/register_d.vhd