../ALU/PFA.vhd