../ALU/barrel_shifter.vhd