../Dataflow/register_file.vhd