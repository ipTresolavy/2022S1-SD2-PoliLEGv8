../Dataflow/mul_div_unit_tb.vhd