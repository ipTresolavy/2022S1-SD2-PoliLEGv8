../Mul_Div_Unit/mul_div_control.vhd