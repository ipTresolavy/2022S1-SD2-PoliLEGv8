../ALU/register_d_bin.vhd