../Dataflow/PFA_tb.vhd