../Dataflow/ALU.vhd