../Mul_Div_Unit/shift_register_tb.vhd