../ALU_pc/ALU_pc.vhd