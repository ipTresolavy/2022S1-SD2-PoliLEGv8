../Dataflow/mux4x1.vhd