../MOV/MOV.vhd