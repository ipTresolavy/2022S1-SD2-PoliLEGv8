../Dataflow/PFA.vhd