../Dataflow/mul_div_unit.vhd