../Dataflow/counter.vhd