../Register_File/register_file.vhd