../Register_File/d_register.vhd