../Dataflow/MOV.vhd