../Dataflow/DataFlow_tb.vhd