../Memory/data_memory_tb.vhd