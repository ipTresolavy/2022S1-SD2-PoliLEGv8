../Dataflow/mux2x1_bin.vhd