../Mul_Div_Unit/mul_div_dataflow.vhd