../Dataflow/barrel_shifter_tb.vhd