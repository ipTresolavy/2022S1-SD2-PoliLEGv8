../ALU/mux2x1.vhd