../Dataflow/data_memory.vhd