../ALU/full_adder.vhd