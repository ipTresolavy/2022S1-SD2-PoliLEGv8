../Memory/instruction_memory.vhd