../Dataflow/ALU_tb.vhd