../Sign_Extension_Unit/sign_extension_unit_tb.vhd