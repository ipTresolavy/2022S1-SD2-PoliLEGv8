../ALU/register_d.vhd