../Dataflow/ALU_4.vhd