../Dataflow/shift_register_tb.vhd