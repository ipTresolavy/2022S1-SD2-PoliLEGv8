../Dataflow/mul_div_control.vhd