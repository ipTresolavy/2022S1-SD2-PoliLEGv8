../Dataflow/DataFlow.vhd