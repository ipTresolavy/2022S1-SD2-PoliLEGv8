../Dataflow/mul_div_dataflow.vhd