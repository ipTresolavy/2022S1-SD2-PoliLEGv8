../Mul_Div_Unit/counter.vhd