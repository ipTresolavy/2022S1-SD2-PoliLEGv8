../Dataflow/register_d_bin.vhd