../Dataflow/mux2x1.vhd