../Mul_Div_Unit/mul_div_unit.vhd